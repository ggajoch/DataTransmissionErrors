library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library unisim;
use unisim.vcomponents.all;

entity clockController is
	port (
		speed_integer : in integer range 10 to 99;
		speed_exp : in integer range 0 to 9;
		clock_100MHz : in std_logic;
		clock_out : out std_logic;
		reset_presc : in std_logic;
		fast_clock : out std_logic
	);
end entity clockController;


architecture RTL of clockController is
	type LUT_Sources_t is array(10 to 729) of integer;
	signal LUT_Sources : LUT_Sources_t := (1, 5, 4, 3, 1, 4, 1, 1, 4, 12, 1, 8, 5, 2, 4, 1, 3, 4, 1, 3, 4, 3, 2, 5, 1, 1, 4, 12, 5, 11, 1, 3, 8, 4, 5, 4, 3, 5, 4, 9, 1, 1, 3, 10, 4, 5, 1, 2, 6, 2, 4, 2, 3, 3, 5, 3, 5, 3, 5, 2, 1, 12, 4, 2, 4, 4, 1, 12, 11, 9, 1, 9, 6, 9, 2, 2, 4, 3, 5, 2, 4, 12, 8, 10, 2, 3, 4, 1, 9, 5, 1, 5, 4, 3, 1, 4, 2, 12, 4, 3, 1, 6, 5, 1, 4, 1, 3, 4, 1, 2, 4, 3, 5, 5, 10, 1, 4, 6, 12, 4, 1, 9, 8, 6, 5, 4, 5, 2, 4, 10, 1, 5, 3, 5, 4, 5, 1, 6, 9, 2, 4, 3, 3, 8, 6, 3, 5, 6, 3, 1, 1, 6, 4, 12, 6, 4, 5, 6, 6, 4, 2, 9, 9, 6, 8, 1, 6, 10, 5, 7, 4, 5, 4, 7, 2, 2, 5, 7, 2, 5, 1, 5, 4, 3, 1, 4, 5, 1, 4, 3, 1, 7, 5, 8, 4, 1, 3, 4, 1, 2, 4, 2, 6, 5, 5, 1, 4, 3, 3, 2, 2, 3, 6, 5, 5, 4, 6, 2, 5, 9, 1, 1, 3, 3, 4, 5, 7, 3, 1, 2, 4, 1, 10, 3, 6, 3, 5, 5, 7, 1, 1, 2, 4, 2, 2, 4, 12, 11, 2, 3, 5, 9, 3, 11, 8, 12, 2, 9, 5, 9, 4, 5, 4, 1, 1, 7, 6, 4, 4, 5, 1, 5, 4, 3, 1, 4, 6, 10, 4, 2, 2, 12, 5, 2, 5, 4, 3, 4, 8, 11, 4, 9, 6, 5, 3, 1, 4, 12, 3, 12, 5, 2, 7, 10, 5, 4, 2, 6, 6, 2, 4, 7, 3, 9, 4, 5, 2, 11, 3, 2, 4, 7, 1, 12, 12, 3, 5, 6, 2, 2, 1, 1, 5, 3, 4, 4, 3, 12, 2, 11, 6, 9, 10, 5, 7, 1, 4, 3, 5, 2, 4, 12, 3, 6, 7, 7, 6, 10, 2, 5, 4, 5, 5, 3, 10, 4, 6, 5, 4, 7, 6, 2, 5, 4, 6, 4, 3, 4, 8, 4, 4, 9, 12, 5, 10, 2, 5, 6, 7, 8, 6, 12, 12, 1, 5, 4, 8, 3, 6, 4, 4, 3, 2, 4, 4, 2, 9, 2, 2, 2, 6, 6, 10, 2, 9, 5, 5, 5, 1, 1, 9, 8, 7, 2, 6, 4, 2, 6, 8, 4, 6, 9, 2, 7, 4, 1, 2, 10, 3, 1, 4, 5, 5, 9, 8, 6, 1, 5, 4, 5, 6, 2, 6, 8, 9, 4, 12, 5, 7, 1, 6, 5, 3, 11, 6, 4, 4, 4, 9, 9, 6, 7, 9, 12, 5, 1, 7, 4, 4, 8, 6, 2, 5, 2, 3, 4, 11, 4, 11, 5, 6, 4, 10, 6, 5, 2, 9, 4, 9, 4, 6, 9, 1, 5, 9, 7, 2, 5, 2, 2, 4, 9, 8, 12, 4, 4, 4, 3, 3, 5, 12, 5, 8, 8, 5, 1, 2, 4, 3, 9, 12, 1, 2, 10, 3, 1, 10, 4, 5, 12, 6, 2, 6, 7, 2, 6, 8, 10, 11, 3, 6, 2, 2, 5, 2, 6, 7, 12, 2, 8, 6, 8, 6, 2, 10, 10, 5, 2, 3, 8, 12, 1, 2, 2, 2, 2, 1, 3, 5, 7, 6, 3, 9, 7, 9, 7, 2, 7, 11, 9, 6, 5, 8, 10, 3, 7, 2, 12, 8, 5, 10, 2, 5, 11, 2, 6, 8, 2, 3, 6, 8, 9, 3, 6, 2, 10, 9, 9, 2, 4, 7, 12, 1, 9, 3, 7, 1, 8, 2, 5, 6, 7, 1, 7, 4, 6, 1, 10, 7, 4, 12, 4, 11, 2, 1, 6, 9, 8, 4, 7, 6, 2, 1, 12, 8, 3, 7, 2, 6, 1, 5, 4, 4, 9, 3, 3, 2, 7, 1, 1, 6, 6, 5, 5, 11, 11, 4, 4, 10, 10, 3, 2, 2, 1, 1, 9, 9, 8, 8, 8, 7, 7, 7, 7, 6, 6, 6, 6, 5, 5, 5, 5, 4, 4, 4, 4, 4, 3, 3, 3, 3, 2, 2, 2, 2, 1, 1, 1, 1, 12);
	



	type LUT_Dividers_t is array(10 to 729) of integer;
	signal LUT_Dividers : LUT_Dividers_t := (192857000, 144360000, 140625000, 137420000, 137755000, 112500000, 120535625, 113445294, 93750000, 52631579, 96428500, 64814762, 72180000, 80393913, 70312500, 77142800, 68710000, 62500000, 68877500, 61602069, 56250000, 57627742, 57783125, 48120000, 56722647, 55102000, 46875000, 27027027, 41788421, 28188718, 48214250, 43572195, 32407381, 39244186, 36090000, 37500000, 38836087, 33786383, 35156250, 26515102, 38571400, 37815098, 34355000, 22471132, 31250000, 28872000, 34438750, 32439649, 25862069, 31340000, 28125000, 30312459, 28813871, 28356508, 24811875, 27484000, 24060000, 26663582, 23352353, 26797971, 27551000, 14084507, 23437500, 25329589, 22804054, 22500000, 25375921, 12987013, 14094359, 16446076, 24107125, 16040000, 18292683, 15653494, 22012619, 21753647, 19622093, 20534023, 18045000, 20775955, 18750000, 10989011, 14794674, 12806129, 19670851, 18804842, 17578125, 19882165, 13257551, 16040000, 19285700, 14436000, 14062500, 13742000, 13775500, 11250000, 11556625, 5882353, 9375000, 9402421, 9642850, 7142857, 7218000, 8385087, 7031250, 7714280, 6871000, 6250000, 6887750, 6376069, 5625000, 5762774, 4962375, 4812000, 3502853, 5510200, 4687500, 4054054, 2631579, 4326923, 4821425, 3168878, 3240738, 3488372, 3609000, 3750000, 3452087, 3934170, 3515625, 2430551, 3857140, 3113647, 3435500, 2996151, 3125000, 2887200, 3443875, 2631579, 2240069, 3134000, 2812500, 2928623, 2881387, 2160492, 2343750, 2748400, 2406000, 2238806, 2627147, 2795029, 2755100, 2112676, 2343750, 1369863, 2027027, 2250000, 2089421, 1948052, 1923077, 2136076, 2311325, 1604000, 1584439, 1807229, 1620369, 2268906, 1744186, 1368931, 1804500, 1605809, 1875000, 1745011, 1834239, 1536742, 1967085, 1946379, 1654125, 1473371, 1886796, 1604000, 1928570, 1443600, 1406250, 1374200, 1377550, 1125000, 992475, 1134453, 937500, 940242, 964285, 680557, 721800, 591787, 703125, 771428, 687100, 625000, 688775, 637607, 562500, 596471, 468750, 481200, 467047, 551020, 468750, 482827, 470121, 474118, 462265, 435722, 357143, 369293, 360900, 375000, 326087, 393417, 330825, 265151, 385714, 378151, 343550, 337068, 312500, 288720, 255209, 313414, 332512, 313400, 281250, 316159, 192092, 283565, 234375, 274840, 240600, 237009, 210172, 279503, 275510, 260431, 234375, 253296, 249873, 225000, 131579, 142774, 237059, 226134, 198495, 160400, 217861, 132453, 162037, 117647, 215007, 149338, 180450, 145982, 187500, 174501, 183424, 207373, 205167, 150439, 156250, 173969, 172194, 160400, 192857, 144360, 140625, 137420, 137755, 112500, 93750, 70057, 93750, 97319, 92453, 47619, 72180, 80394, 66165, 67500, 68710, 62500, 48611, 37909, 56250, 41911, 46875, 48120, 52543, 55102, 46875, 27027, 47012, 25641, 39699, 45099, 34028, 27697, 36090, 37500, 40197, 31915, 31250, 37736, 33750, 28023, 34355, 24514, 31250, 28872, 33019, 19287, 30801, 31340, 28125, 23429, 31106, 15873, 15625, 27484, 24060, 22388, 27192, 26798, 27551, 27163, 22055, 24472, 22804, 22500, 23506, 12987, 23706, 13916, 18750, 16040, 14524, 19132, 17014, 22689, 19622, 20534, 18045, 20776, 18750, 10989, 19418, 16129, 15204, 15044, 15625, 12278, 18868, 16040, 16875, 14436, 13233, 13742, 8507, 11250, 9375, 9341, 9375, 7522, 7500, 8805, 7218, 7337, 6250, 6750, 6871, 6250, 4861, 5819, 5625, 4191, 3125, 4812, 3503, 5283, 4411, 4054, 3761, 3490, 3750, 2439, 2381, 4485, 3609, 3750, 2959, 3801, 3125, 3444, 3375, 3503, 3556, 3184, 3125, 3362, 2320, 3244, 3188, 3134, 2500, 2459, 1921, 2935, 2030, 2443, 2406, 2370, 2836, 2795, 1856, 1917, 1985, 2533, 2027, 2250, 2433, 1948, 1745, 2136, 1875, 1604, 2255, 1722, 2009, 2269, 2150, 1369, 2030, 2167, 1875, 1745, 1726, 1397, 1448, 1579, 2009, 1637, 1722, 1604, 1500, 1681, 1250, 1047, 928, 1125, 625, 934, 794, 1015, 750, 756, 812, 478, 625, 675, 649, 625, 464, 448, 500, 461, 406, 303, 467, 551, 397, 456, 444, 349, 375, 451, 378, 430, 406, 375, 239, 359, 229, 324, 300, 331, 229, 283, 294, 336, 232, 296, 224, 286, 250, 213, 311, 252, 203, 220, 280, 237, 272, 268, 241, 183, 189, 137, 228, 225, 222, 232, 229, 201, 125, 196, 166, 164, 189, 227, 215, 194, 203, 146, 111, 212, 201, 128, 190, 203, 124, 174, 162, 101, 150, 168, 125, 110, 132, 100, 85, 70, 61, 94, 75, 88, 84, 69, 77, 60, 55, 37, 66, 47, 50, 44, 47, 56, 35, 34, 44, 50, 47, 35, 25, 47, 44, 43, 42, 41, 42, 38, 33, 29, 30, 35, 25, 27, 24, 26, 33, 25, 19, 22, 25, 26, 22, 19, 28, 22, 28, 15, 20, 23, 17, 26, 22, 15, 25, 20, 18, 24, 23, 19, 17, 16, 22, 18, 22, 14, 15, 15, 21, 19, 16, 11, 21, 14, 19, 15, 20, 14, 19, 16, 15, 13, 16, 11, 12, 10, 12, 7, 8, 9, 5, 8, 5, 8, 8, 6, 5, 5, 6, 5, 5, 6, 6, 3, 4, 5, 4, 5, 4, 5, 4, 4, 4, 3, 4, 4, 4, 3, 4, 4, 3, 3, 3, 3, 2, 2, 3, 3, 2, 2, 3, 3, 3, 3, 3, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 1);




	
	
	--400e6, 390e6, 360e6, 350e6, 340e6, 320e6, 300e6, 250e6
	signal PLL_vals : std_logic_vector(1 to 13);
	
	signal presc_in : std_logic;
	signal presc_in_unbuffered : std_logic;
	signal presc_out : std_logic;
	signal presc_rst : std_logic;
	signal presc_val : integer;
	signal index : integer range 10 to 730;
	
	component clk_wiz_0
    port
     (-- Clock in ports
      clk_in1           : in     std_logic;
      -- Clock out ports
      clk_out1          : out    std_logic;
      clk_out2          : out    std_logic;
      clk_out3          : out    std_logic;
      clk_out4          : out    std_logic;
      clk_out5          : out    std_logic;
      clk_out6          : out    std_logic
     );
    end component;
    
    ATTRIBUTE SYN_BLACK_BOX : BOOLEAN;
    ATTRIBUTE SYN_BLACK_BOX OF clk_wiz_0 : COMPONENT IS TRUE;
    ATTRIBUTE BLACK_BOX_PAD_PIN : STRING;
    ATTRIBUTE BLACK_BOX_PAD_PIN OF clk_wiz_0 : COMPONENT IS "clk_in1,clk_out1,clk_out2,clk_out3,clk_out4,clk_out5,clk_out6";
    
    
    component clk_wiz_1
    port
     (-- Clock in ports
      clk_in1           : in     std_logic;
      -- Clock out ports
      clk_out1          : out    std_logic;
      clk_out2          : out    std_logic;
      clk_out3          : out    std_logic
     );
    end component;
    
    --ATTRIBUTE SYN_BLACK_BOX : BOOLEAN;
    ATTRIBUTE SYN_BLACK_BOX OF clk_wiz_1 : COMPONENT IS TRUE;
    --ATTRIBUTE BLACK_BOX_PAD_PIN : STRING;
    ATTRIBUTE BLACK_BOX_PAD_PIN OF clk_wiz_1 : COMPONENT IS "clk_in1,clk_out1,clk_out2,clk_out3";
    
    
    
    component clk_wiz_2
    port
     (-- Clock in ports
      clk_in1           : in     std_logic;
      -- Clock out ports
      clk_out1          : out    std_logic;
      clk_out2          : out    std_logic
     );
    end component;
    
    --ATTRIBUTE SYN_BLACK_BOX : BOOLEAN;
    ATTRIBUTE SYN_BLACK_BOX OF clk_wiz_2 : COMPONENT IS TRUE;
    --ATTRIBUTE BLACK_BOX_PAD_PIN : STRING;
    ATTRIBUTE BLACK_BOX_PAD_PIN OF clk_wiz_2 : COMPONENT IS "clk_in1,clk_out1,clk_out2";

begin
	
	--------------- PLL -----------------
	
	--PLL_vals <= clock_100MHz & clock_100MHz & clock_100MHz & clock_100MHz & clock_100MHz & clock_100MHz & clock_100MHz & clock_100MHz;
	
	PLL0_inst : clk_wiz_0
       port map ( 
    
       -- Clock in ports
       clk_in1 => clock_100MHz,
      -- Clock out ports  
       clk_out1 => PLL_vals(11),
       clk_out2 => PLL_vals(10),
       clk_out3 => PLL_vals(9),
       clk_out4 => PLL_vals(7),
       clk_out5 => PLL_vals(5),
       clk_out6 => PLL_vals(3)              
     );
     
     PLL1_inst : clk_wiz_1
        port map ( 
     
        -- Clock in ports
        clk_in1 => clock_100MHz,
       -- Clock out ports  
        clk_out1 => PLL_vals(6),
        clk_out2 => PLL_vals(4),
        clk_out3 => PLL_vals(1)
      );
      
      PLL2_inst : clk_wiz_2
          port map ( 
       
          -- Clock in ports
          clk_in1 => clock_100MHz,
         -- Clock out ports  
          clk_out1 => PLL_vals(2),
          clk_out2 => PLL_vals(8)             
        );
	
	PLL_vals(12) <= clock_100MHz;
	------------- PRESCALER -------------
	
	fast_clock <= PLL_vals(9);
	
	index <= speed_integer + 90*speed_exp;
	presc_in_unbuffered <= PLL_vals(LUT_Sources(index));
	presc_val <= LUT_Dividers(index);

	presc_rst <= reset_presc;
	
	presc_in_buf : BUFG
               port map
                (O   => presc_in,
                 I   => presc_in_unbuffered);
	
	presc_inst : entity work.prescaler
		port map(clk_input  => presc_in,
			     clk_output => presc_out,
			     reset      => presc_rst,
			     presc      => presc_val);
	
	
	
	------------- BUFG -----------------
	--clock_out <= presc_out;
	
	clkout1_buf : BUFG
           port map
            (O   => clock_out,
             I   => presc_out);

end architecture RTL;
