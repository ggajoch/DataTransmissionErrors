library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library unisim;
use unisim.vcomponents.all;

entity clockController is
	port (
		speed_integer : in integer range 10 to 99;
		speed_exp : in integer range 0 to 9;
		clock_100MHz : in std_logic;
		clock_out : out std_logic;
		reset_presc : in std_logic;
		fast_clock : out std_logic
	);
end entity clockController;


architecture RTL of clockController is
	type LUT_Sources_t is array(10 to 729) of integer;
	signal LUT_Sources : LUT_Sources_t := (1, 1, 1, 2, 4, 1, 1, 4, 1, 6, 1, 6, 1, 3, 1, 1, 2, 6, 4, 1, 1, 2, 4, 1, 4, 4, 1, 4, 1, 2, 1, 4, 6, 6, 1, 1, 4, 2, 1, 5, 1, 2, 2, 6, 6, 1, 4, 6, 1, 5, 1, 1, 4, 6, 1, 2, 1, 3, 4, 3, 4, 3, 1, 1, 4, 1, 3, 3, 2, 1, 1, 5, 2, 2, 1, 4, 1, 1, 1, 1, 1, 1, 2, 4, 2, 5, 3, 3, 3, 1, 1, 1, 1, 2, 4, 1, 4, 4, 1, 3, 1, 5, 1, 2, 1, 1, 2, 2, 4, 1, 1, 1, 1, 1, 4, 4, 1, 4, 6, 2, 1, 5, 6, 5, 1, 1, 1, 4, 3, 3, 1, 2, 2, 4, 2, 1, 4, 4, 1, 4, 1, 2, 1, 2, 3, 2, 1, 3, 4, 3, 4, 4, 1, 1, 4, 1, 1, 2, 2, 4, 4, 2, 5, 3, 6, 4, 4, 1, 1, 2, 1, 4, 1, 4, 2, 2, 3, 2, 1, 1, 1, 1, 1, 2, 4, 1, 1, 4, 1, 5, 1, 3, 1, 3, 3, 1, 2, 3, 4, 1, 1, 1, 1, 1, 4, 4, 1, 4, 3, 2, 4, 1, 5, 6, 1, 1, 4, 6, 6, 3, 1, 1, 2, 3, 4, 1, 4, 5, 1, 3, 1, 6, 1, 3, 5, 2, 1, 3, 4, 2, 4, 2, 2, 1, 4, 1, 6, 3, 2, 1, 1, 3, 1, 4, 6, 4, 5, 1, 4, 6, 1, 1, 2, 1, 6, 4, 5, 1, 4, 1, 1, 1, 3, 2, 4, 1, 3, 4, 1, 2, 4, 3, 1, 1, 3, 6, 2, 6, 4, 1, 1, 4, 3, 1, 4, 4, 6, 4, 5, 2, 1, 1, 3, 3, 3, 1, 3, 2, 3, 1, 6, 1, 3, 1, 6, 1, 3, 1, 1, 3, 3, 1, 3, 5, 6, 2, 1, 1, 4, 3, 4, 3, 4, 1, 4, 3, 2, 3, 2, 5, 1, 3, 1, 1, 3, 4, 6, 1, 3, 5, 1, 1, 3, 4, 1, 4, 3, 2, 1, 1, 5, 1, 6, 2, 4, 4, 1, 4, 3, 4, 2, 1, 5, 4, 5, 4, 1, 2, 1, 1, 4, 3, 3, 1, 4, 1, 1, 4, 6, 2, 2, 2, 1, 1, 5, 5, 1, 3, 5, 4, 4, 6, 5, 6, 1, 6, 5, 1, 4, 1, 4, 2, 3, 1, 3, 3, 2, 1, 2, 3, 1, 2, 1, 1, 4, 4, 6, 2, 1, 1, 2, 2, 3, 2, 1, 5, 1, 1, 4, 4, 2, 4, 1, 3, 3, 1, 1, 2, 6, 1, 4, 4, 2, 1, 1, 4, 1, 1, 2, 1, 5, 1, 3, 4, 1, 5, 1, 2, 5, 4, 4, 1, 1, 5, 3, 3, 1, 3, 2, 2, 1, 3, 1, 4, 3, 3, 2, 1, 5, 2, 5, 1, 1, 2, 2, 1, 5, 2, 4, 3, 2, 6, 1, 5, 3, 2, 4, 2, 3, 4, 4, 3, 1, 2, 3, 2, 4, 1, 2, 3, 1, 1, 3, 2, 5, 6, 4, 4, 4, 2, 3, 5, 2, 4, 1, 5, 3, 2, 2, 2, 5, 4, 6, 2, 4, 2, 1, 4, 3, 5, 1, 2, 4, 5, 2, 2, 2, 6, 1, 2, 2, 2, 2, 2, 4, 3, 2, 3, 3, 2, 6, 5, 1, 6, 4, 5, 3, 3, 4, 2, 2, 1, 4, 3, 2, 1, 2, 5, 1, 2, 1, 2, 1, 2, 1, 2, 5, 3, 4, 5, 3, 4, 2, 5, 4, 2, 3, 5, 2, 4, 1, 2, 5, 4, 1, 2, 2, 1, 4, 2, 6, 1, 3, 2, 5, 1, 1, 6, 2, 4, 1, 1, 5, 2, 1, 2, 1, 6, 2, 1, 2, 1, 5, 1, 2, 3, 1, 5, 2, 6, 1, 1, 2, 5, 1, 3, 3, 4, 4, 2, 2, 1, 1, 3, 5, 5, 5, 2, 2, 2, 4, 4, 1, 1, 1, 1, 6, 6, 6, 3, 3, 3, 2, 2, 2, 2, 5, 5, 1, 1, 1, 1, 1, 4, 4, 4, 4, 4, 4, 4, 4, 4, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 2, 2, 2, 2, 2, 2, 2);



	type LUT_Dividers_t is array(10 to 729) of integer;
	signal LUT_Dividers : LUT_Dividers_t := (209583000, 190530000, 174652500, 149970000, 106930000, 139722000, 130989375, 88060000, 116435000, 61281579, 104791500, 55445238, 95265000, 75936087, 87326250, 83833200, 74985000, 43124074, 53465000, 72270000, 69861000, 62890645, 46781875, 63510000, 44030000, 42772000, 58217500, 40460000, 55153421, 49990000, 52395750, 36512683, 27722619, 27077907, 47632500, 46574000, 32543913, 41481064, 43663125, 26732653, 41916600, 38227647, 37492500, 21968868, 21562037, 38106000, 26732500, 20427193, 36135000, 22201695, 34930500, 34357869, 24145484, 18481746, 32747344, 29994000, 31755000, 26067612, 22015000, 25312029, 21386000, 24599014, 29108750, 28710000, 20230000, 27944400, 22980658, 22682208, 24995000, 26529494, 26197875, 16171605, 23775732, 23489277, 24950357, 17612000, 24370116, 24090000, 23816250, 23548652, 23287000, 23031099, 21191413, 16096989, 20740532, 13788421, 18193021, 18005464, 17821735, 21170000, 20958300, 19053000, 17465250, 14997000, 10693000, 13972200, 9356375, 8806000, 11643500, 9192263, 10479150, 6237619, 9526500, 8476565, 8732625, 8383320, 7498500, 7220778, 5346500, 7227000, 6986100, 6760742, 6549469, 6351000, 4403000, 4277200, 5821750, 4046000, 3064079, 4999000, 5239575, 3194878, 2772262, 3046279, 4763250, 4657400, 4556152, 3185149, 3638604, 3564347, 4191660, 3822765, 3749250, 2824566, 3610389, 3810600, 2673250, 2626351, 3613500, 2537322, 3493050, 3196082, 3380371, 3094619, 2728953, 2999400, 3175500, 2606761, 2201500, 2531203, 2138600, 2108479, 2910875, 2871000, 2023000, 2794440, 2757671, 2531961, 2499500, 1894962, 1871275, 2406926, 1597439, 2104253, 1386131, 1761200, 1740721, 2409000, 2381625, 2190573, 2328700, 1645077, 2278076, 1609699, 2074053, 2052221, 1819302, 2009907, 2138602, 2117000, 2095830, 1905300, 1746525, 1499700, 1069300, 1397220, 1309894, 880600, 1164350, 689421, 1047915, 831681, 952650, 759361, 727721, 838332, 749850, 646863, 534650, 722700, 698610, 676074, 654947, 635100, 440300, 427720, 582175, 404600, 459613, 499900, 374255, 511178, 311881, 270779, 476325, 465740, 325439, 247734, 242573, 356435, 419166, 410947, 374925, 329534, 277226, 381060, 267325, 229807, 361350, 296022, 349305, 190877, 338037, 277227, 204672, 299940, 317550, 260676, 220150, 282552, 213860, 274593, 270779, 287100, 202300, 279444, 153204, 226822, 249950, 265295, 261979, 215621, 255589, 180364, 138613, 176120, 152314, 240900, 170116, 130826, 232870, 230311, 211914, 225358, 123867, 157581, 136448, 216065, 152757, 211700, 209583, 190530, 145544, 149970, 106930, 139722, 109158, 88060, 116435, 102611, 74851, 83168, 95265, 91123, 72772, 46574, 74985, 43124, 53465, 72270, 69861, 48291, 54579, 63510, 44030, 42772, 32343, 40460, 34471, 49990, 52396, 51118, 41584, 40617, 39694, 46574, 37968, 41481, 36386, 42772, 23287, 41095, 33587, 39544, 21562, 38106, 31188, 36769, 36135, 29602, 29109, 34358, 28170, 20792, 18193, 29994, 31755, 31281, 22015, 25312, 21386, 24599, 20792, 28710, 20230, 23287, 25653, 22682, 24995, 16581, 26198, 21562, 25559, 25251, 20792, 17612, 13539, 24090, 19847, 14718, 23287, 23031, 18984, 16097, 22296, 15758, 18193, 20099, 21386, 21170, 13099, 19053, 9703, 14997, 10693, 9980, 13099, 8806, 9703, 7879, 9748, 9980, 5954, 6509, 5458, 5988, 8061, 7221, 7485, 7227, 4990, 5634, 5458, 6351, 4403, 5988, 5822, 4046, 3064, 4999, 4874, 4755, 4990, 4874, 2977, 2911, 4556, 3716, 2729, 3055, 2994, 2283, 2519, 2197, 3881, 2117, 2339, 3677, 2581, 3552, 2495, 3196, 2817, 3327, 2729, 2687, 2954, 3128, 2867, 2531, 2994, 2746, 2911, 2871, 2023, 1996, 1532, 2532, 2687, 2653, 2437, 2407, 2130, 2349, 2495, 1541, 2437, 2409, 1701, 1682, 2166, 1645, 2278, 1878, 1858, 2206, 2183, 2010, 1188, 2117, 1497, 1361, 1625, 1612, 1497, 998, 1310, 1233, 1083, 1103, 655, 998, 794, 651, 873, 524, 806, 722, 468, 516, 499, 676, 655, 397, 514, 499, 582, 472, 513, 500, 524, 426, 499, 348, 397, 388, 424, 446, 273, 398, 262, 411, 403, 368, 361, 381, 234, 342, 258, 296, 325, 191, 338, 208, 273, 300, 227, 291, 257, 217, 214, 246, 291, 267, 236, 260, 197, 272, 250, 221, 262, 259, 213, 235, 156, 137, 174, 172, 170, 219, 194, 144, 212, 161, 223, 138, 182, 201, 199, 197, 131, 136, 97, 150, 107, 130, 131, 88, 97, 69, 105, 93, 68, 57, 81, 78, 75, 43, 75, 67, 65, 63, 61, 59, 44, 50, 54, 47, 46, 50, 29, 32, 50, 27, 34, 29, 38, 37, 31, 40, 39, 41, 29, 33, 36, 38, 35, 23, 36, 33, 35, 32, 34, 31, 33, 30, 20, 26, 22, 19, 25, 21, 27, 18, 20, 26, 23, 17, 25, 19, 26, 24, 16, 18, 25, 23, 23, 24, 17, 22, 13, 23, 19, 21, 14, 22, 22, 12, 20, 15, 21, 19, 11, 15, 15, 13, 13, 7, 11, 11, 10, 10, 6, 9, 8, 7, 8, 5, 7, 4, 7, 7, 6, 4, 6, 5, 5, 4, 4, 5, 5, 5, 5, 4, 3, 3, 3, 4, 4, 4, 3, 3, 4, 4, 4, 4, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 2, 2, 3, 3, 3, 3, 3, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2);



	
	
	--400e6, 390e6, 360e6, 350e6, 340e6, 320e6, 300e6, 250e6
	signal PLL_vals : std_logic_vector(1 to 8);
	
	signal presc_in : std_logic;
	signal presc_in_unbuffered : std_logic;
	signal presc_out : std_logic;
	signal presc_rst : std_logic;
	signal presc_val : integer;
	signal index : integer range 10 to 730;
	
	
	component clk_wiz_0
    port
     (-- Clock in ports
      clk_in1           : in     std_logic;
      -- Clock out ports
      clk_out1          : out    std_logic;
      clk_out2          : out    std_logic;
      clk_out3          : out    std_logic;
      clk_out4          : out    std_logic;
      clk_out5          : out    std_logic;
      clk_out6          : out    std_logic
     );
    end component;
    
    ATTRIBUTE SYN_BLACK_BOX : BOOLEAN;
    ATTRIBUTE SYN_BLACK_BOX OF clk_wiz_0 : COMPONENT IS TRUE;
    
    
    ATTRIBUTE BLACK_BOX_PAD_PIN : STRING;
    ATTRIBUTE BLACK_BOX_PAD_PIN OF clk_wiz_0 : COMPONENT IS "clk_in1,clk_out1,clk_out2,clk_out3,clk_out4,clk_out5,clk_out6";

begin
	
	--------------- PLL -----------------
	
	--PLL_vals <= clock_100MHz & clock_100MHz & clock_100MHz & clock_100MHz & clock_100MHz & clock_100MHz & clock_100MHz & clock_100MHz;
	
	PLL0_inst : clk_wiz_0
       port map ( 
    
       -- Clock in ports
       clk_in1 => clock_100MHz,
      -- Clock out ports  
       clk_out1 => PLL_vals(1),
       clk_out2 => PLL_vals(2),
       clk_out3 => PLL_vals(3),
       clk_out4 => PLL_vals(4),
       clk_out5 => PLL_vals(5),
       clk_out6 => PLL_vals(6)              
     );
	
	------------- PRESCALER -------------
	
	fast_clock <= PLL_vals(1);
	
	index <= speed_integer + 90*speed_exp;
	presc_in_unbuffered <= PLL_vals(LUT_Sources(index));
	presc_val <= LUT_Dividers(index);

	presc_rst <= reset_presc;
	
	presc_in_buf : BUFG
               port map
                (O   => presc_in,
                 I   => presc_in_unbuffered);
	
	presc_inst : entity work.prescaler
		port map(clk_input  => presc_in,
			     clk_output => presc_out,
			     reset      => presc_rst,
			     presc      => presc_val);
	
	
	
	------------- BUFG -----------------
	--clock_out <= presc_out;
	
	clkout1_buf : BUFG
           port map
            (O   => clock_out,
             I   => presc_out);

end architecture RTL;
