library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library unisim;
use unisim.vcomponents.all;

entity clockController is
	port (
		speed_integer : in integer range 10 to 99;
		speed_exp : in integer range 0 to 9;
		clock_100MHz : in std_logic;
		clock_out : out std_logic;
		reset_presc : in std_logic
	);
end entity clockController;


architecture RTL of clockController is
	type LUT_Sources_t is array(10 to 729) of integer;
    signal LUT_Sources : LUT_Sources_t := (1, 2, 1, 2, 1, 1, 1, 6, 3, 6, 1, 1, 2, 2, 1, 1, 2, 7, 1, 4, 1, 4, 1, 4, 4, 1, 3, 2, 6, 3, 1, 4, 1, 1, 2, 3, 2, 2, 1, 6, 1, 6, 2, 7, 7, 2, 1, 6, 4, 1, 1, 6, 4, 3, 2, 2, 4, 7, 4, 5, 1, 7, 3, 6, 2, 1, 1, 2, 3, 7, 1, 1, 4, 1, 1, 1, 6, 2, 2, 4, 3, 2, 1, 1, 1, 3, 1, 2, 6, 5, 1, 2, 1, 2, 1, 1, 1, 2, 3, 3, 1, 1, 2, 3, 1, 1, 2, 7, 1, 1, 1, 5, 2, 4, 2, 1, 3, 2, 6, 3, 1, 2, 1, 1, 2, 3, 7, 7, 1, 6, 1, 4, 2, 4, 7, 2, 1, 1, 3, 2, 1, 1, 5, 3, 6, 2, 4, 1, 2, 1, 1, 1, 3, 1, 2, 1, 6, 2, 3, 6, 1, 5, 2, 1, 1, 6, 5, 4, 2, 7, 3, 2, 1, 5, 4, 3, 3, 2, 6, 7, 1, 2, 1, 2, 1, 1, 2, 4, 3, 3, 1, 1, 2, 2, 1, 1, 2, 7, 1, 7, 1, 2, 6, 4, 4, 1, 3, 2, 3, 3, 1, 1, 1, 2, 2, 3, 2, 5, 3, 6, 1, 7, 2, 3, 7, 2, 1, 1, 5, 5, 1, 7, 5, 3, 6, 2, 4, 6, 1, 2, 1, 2, 3, 1, 2, 1, 6, 2, 3, 3, 2, 4, 2, 1, 1, 2, 2, 1, 2, 1, 3, 2, 3, 2, 3, 4, 7, 2, 6, 5, 1, 2, 1, 2, 1, 1, 6, 2, 3, 3, 1, 1, 2, 1, 3, 1, 2, 7, 1, 4, 1, 1, 6, 4, 2, 1, 3, 2, 3, 3, 2, 1, 1, 2, 2, 3, 2, 2, 7, 6, 1, 1, 2, 1, 7, 2, 2, 2, 4, 1, 1, 4, 1, 3, 6, 2, 4, 1, 4, 3, 1, 2, 3, 5, 2, 1, 3, 2, 3, 2, 6, 6, 1, 1, 1, 4, 4, 7, 2, 6, 3, 2, 2, 2, 3, 4, 2, 2, 6, 7, 1, 2, 3, 2, 1, 1, 6, 4, 3, 4, 5, 1, 2, 3, 7, 5, 2, 7, 2, 1, 1, 2, 6, 4, 4, 1, 3, 2, 4, 3, 6, 4, 1, 4, 2, 7, 3, 3, 1, 6, 5, 2, 2, 3, 7, 1, 6, 2, 1, 2, 7, 3, 3, 3, 6, 7, 5, 1, 4, 2, 1, 4, 7, 6, 2, 7, 4, 2, 3, 1, 6, 2, 4, 2, 3, 3, 4, 2, 6, 3, 7, 2, 7, 2, 2, 1, 1, 2, 6, 5, 5, 3, 7, 7, 5, 7, 6, 3, 7, 3, 6, 1, 3, 3, 4, 1, 7, 7, 6, 3, 7, 3, 6, 2, 1, 5, 7, 1, 3, 7, 6, 4, 2, 1, 5, 7, 1, 3, 1, 6, 1, 4, 7, 6, 7, 4, 6, 5, 3, 7, 7, 2, 2, 2, 5, 7, 1, 6, 1, 1, 5, 1, 6, 3, 6, 1, 5, 1, 7, 1, 6, 2, 1, 3, 1, 1, 3, 1, 5, 1, 7, 4, 1, 1, 3, 2, 7, 3, 6, 7, 2, 4, 3, 7, 6, 1, 6, 1, 7, 2, 2, 4, 3, 1, 5, 1, 7, 7, 6, 6, 4, 3, 7, 5, 1, 7, 1, 2, 2, 7, 2, 2, 3, 4, 7, 2, 6, 7, 2, 6, 1, 2, 6, 2, 7, 3, 6, 2, 3, 2, 6, 3, 2, 1, 7, 6, 1, 2, 1, 4, 7, 6, 3, 1, 2, 3, 1, 1, 7, 1, 4, 5, 2, 1, 1, 4, 4, 6, 7, 5, 1, 1, 2, 3, 3, 1, 1, 6, 6, 5, 1, 3, 1, 6, 7, 3, 4, 1, 5, 1, 3, 1, 4, 7, 1, 2, 6, 1, 4, 2, 3, 3, 1, 1, 7, 7, 7, 2, 1, 6, 3, 3, 3, 5, 5, 5, 5, 1, 1, 2, 2, 2, 2, 4, 4, 4, 4, 4, 4, 3, 3, 3, 3, 1, 1, 1, 1, 7, 7, 7, 7, 7, 7, 2, 2, 2, 2, 6, 6, 6, 6, 6, 6, 6, 5, 5, 5, 5, 5, 5, 5, 5, 5, 1, 1, 1, 1, 1, 1, 1);

	type LUT_Dividers_t is array(10 to 729) of integer;
    signal LUT_Dividers : LUT_Dividers_t := (190470000, 134680000, 158725000, 113960000, 136050000, 126980000, 119043750, 46117647, 67340000, 41263158, 95235000, 90700000, 67340000, 64412174, 79362500, 76188000, 56980000, 26000000, 68025000, 38314138, 63490000, 35842258, 59521875, 33670000, 32679706, 54420000, 33670000, 40040000, 20631579, 31080000, 47617500, 27100244, 45350000, 44295349, 33670000, 26936000, 32206087, 31520851, 39681250, 16000000, 38094000, 15372549, 28490000, 13245283, 13000000, 26936000, 34012500, 13754386, 19157069, 32283051, 31745000, 12852459, 17921129, 19240000, 23148125, 22792000, 16835000, 10477612, 16339853, 12884058, 27210000, 9887324, 16835000, 10739726, 20020000, 25396000, 25061842, 19240000, 15540000, 8886076, 23808750, 23514815, 13550122, 22948193, 22675000, 22408235, 9116279, 17028506, 16835000, 12484382, 13468000, 16280000, 20703261, 20480645, 20262766, 12759158, 19840625, 15272990, 8000000, 8979798, 19047000, 13468000, 15872500, 11396000, 13605000, 12698000, 11904375, 8714588, 6734000, 6379579, 9523500, 9070000, 6734000, 5270087, 7936250, 7618800, 5698000, 2600000, 6802500, 6567931, 6349000, 2867742, 4629625, 3367000, 4357294, 5442000, 3367000, 4004000, 2063158, 3108000, 4761750, 3613366, 4535000, 4429535, 3367000, 2693600, 1526087, 1493617, 3968125, 1600000, 3809400, 2178647, 2849000, 2096434, 1300000, 2693600, 3401250, 3341579, 2089862, 2510983, 3174500, 3122459, 1433871, 1924000, 1225000, 2279200, 1683500, 2842836, 2178647, 2760435, 2721000, 2682676, 1683500, 2609178, 2002000, 2539600, 1031579, 1924000, 1554000, 992405, 2380875, 1097531, 1806683, 2294819, 2267500, 922353, 1033721, 1277138, 1683500, 788764, 1346800, 1628000, 2070326, 955914, 1182032, 1275916, 1262625, 1527299, 800000, 709091, 1904700, 1346800, 1587250, 1139600, 1360500, 1269800, 925925, 653594, 673400, 637958, 952350, 907000, 673400, 644122, 793625, 761880, 569800, 260000, 680250, 242069, 634900, 477897, 245000, 336700, 326797, 544200, 336700, 400400, 318979, 310800, 476175, 464561, 453500, 344530, 336700, 269360, 322061, 189149, 252525, 160000, 380940, 137647, 284900, 228702, 130000, 269360, 340125, 334158, 153276, 150678, 317450, 115082, 143387, 192400, 122500, 227920, 168350, 117015, 280103, 214707, 272100, 208659, 168350, 260918, 200200, 253960, 103158, 192400, 155400, 153433, 185185, 137174, 180668, 229482, 226750, 174292, 172265, 218931, 168350, 214011, 134680, 162800, 131752, 159299, 128949, 116959, 73125, 152730, 80000, 89798, 190470, 134680, 158725, 113960, 136050, 126980, 49000, 87146, 67340, 63796, 95235, 90700, 67340, 82813, 50505, 76188, 56980, 26000, 68025, 38314, 63490, 61442, 24500, 33670, 43573, 54420, 33670, 40040, 31898, 31080, 37037, 46456, 45350, 34453, 33670, 26936, 32206, 31521, 14625, 16000, 38094, 37347, 28490, 35938, 13000, 26936, 26455, 25991, 19157, 32283, 31745, 18215, 30721, 19240, 12250, 22792, 16835, 28428, 16340, 17567, 27210, 20866, 16835, 12178, 20020, 25396, 15949, 19240, 15540, 18753, 9800, 9679, 23228, 22948, 22675, 13072, 12920, 8069, 16835, 8809, 13468, 16280, 16103, 15930, 12895, 11696, 15432, 15273, 8000, 7091, 19047, 13468, 10101, 11396, 13605, 12698, 4900, 6536, 6734, 5848, 4445, 9070, 6734, 5270, 2925, 3556, 5698, 2600, 5291, 6568, 6349, 4779, 2450, 3367, 3268, 5442, 3367, 4004, 2924, 3108, 1960, 2710, 4535, 2584, 3367, 1560, 2635, 2579, 3968, 1600, 1778, 2905, 2849, 2287, 1300, 3463, 1400, 2599, 3284, 2511, 1170, 1987, 1955, 1924, 1225, 1080, 1347, 2843, 1634, 2147, 2721, 1565, 975, 1074, 2002, 936, 1462, 1924, 1554, 2411, 980, 1829, 1355, 1785, 1443, 1426, 1292, 1703, 891, 1362, 780, 1628, 763, 1593, 1576, 2005, 1984, 1527, 800, 898, 889, 1102, 585, 540, 635, 468, 490, 713, 390, 638, 392, 907, 551, 527, 463, 762, 270, 260, 280, 418, 234, 391, 245, 449, 560, 254, 195, 515, 319, 180, 196, 271, 353, 443, 202, 156, 414, 258, 397, 160, 381, 218, 135, 148, 130, 202, 140, 156, 209, 119, 117, 243, 239, 235, 139, 108, 289, 117, 280, 276, 127, 268, 109, 166, 106, 254, 117, 247, 90, 241, 98, 183, 232, 146, 227, 224, 141, 219, 101, 214, 78, 122, 207, 205, 129, 156, 73, 125, 80, 71, 148, 101, 101, 54, 56, 127, 49, 112, 39, 78, 74, 53, 55, 83, 37, 76, 27, 26, 28, 27, 37, 39, 22, 27, 56, 20, 53, 40, 39, 18, 37, 36, 29, 26, 16, 33, 17, 15, 31, 16, 38, 29, 15, 28, 13, 22, 14, 26, 21, 25, 13, 20, 24, 30, 11, 12, 29, 22, 28, 16, 10, 11, 17, 26, 20, 16, 25, 25, 9, 24, 14, 11, 18, 23, 23, 13, 13, 9, 8, 10, 21, 21, 16, 13, 13, 20, 20, 8, 8, 9, 19, 11, 16, 6, 5, 8, 7, 11, 5, 10, 6, 9, 5, 3, 8, 6, 3, 7, 4, 5, 4, 4, 6, 6, 2, 2, 2, 4, 5, 2, 3, 3, 3, 2, 2, 2, 2, 4, 4, 3, 3, 3, 3, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 3, 3, 3, 3, 1, 1, 1, 1, 1, 1, 2, 2, 2, 2, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2);

	
	
	--400e6, 390e6, 360e6, 350e6, 340e6, 320e6, 300e6, 250e6
	signal PLL_vals : std_logic_vector(1 to 8);
	
	signal presc_in : std_logic;
	signal presc_in_unbuffered : std_logic;
	signal presc_out : std_logic;
	signal presc_rst : std_logic;
	signal presc_val : integer;
	signal index : integer range 10 to 730;
	
	
	component clk_wiz_0
    port
     (-- Clock in ports
      clk_in1           : in     std_logic;
      -- Clock out ports
      clk_out1          : out    std_logic;
      clk_out2          : out    std_logic;
      clk_out3          : out    std_logic;
      clk_out4          : out    std_logic;
      clk_out5          : out    std_logic;
      clk_out6          : out    std_logic;
      clk_out7          : out    std_logic
     );
    end component;
    
    ATTRIBUTE SYN_BLACK_BOX : BOOLEAN;
    ATTRIBUTE SYN_BLACK_BOX OF clk_wiz_0 : COMPONENT IS TRUE;
    
    
    ATTRIBUTE BLACK_BOX_PAD_PIN : STRING;
    ATTRIBUTE BLACK_BOX_PAD_PIN OF clk_wiz_0 : COMPONENT IS "clk_in1,clk_out1,clk_out2,clk_out3,clk_out4,clk_out5,clk_out6,clk_out7";

begin
	
	--------------- PLL -----------------
	
	--PLL_vals <= clock_100MHz & clock_100MHz & clock_100MHz & clock_100MHz & clock_100MHz & clock_100MHz & clock_100MHz & clock_100MHz;
	
	PLL0_inst : clk_wiz_0
       port map ( 
    
       -- Clock in ports
       clk_in1 => clock_100MHz,
      -- Clock out ports  
       clk_out1 => PLL_vals(1),
       clk_out2 => PLL_vals(2),
       clk_out3 => PLL_vals(3),
       clk_out4 => PLL_vals(4),
       clk_out5 => PLL_vals(5),
       clk_out6 => PLL_vals(6),
       clk_out7 => PLL_vals(7)              
     );
	
	------------- PRESCALER -------------
	
	index <= speed_integer + 90*speed_exp;
	presc_in_unbuffered <= PLL_vals(LUT_Sources(index));
	presc_val <= LUT_Dividers(index);

	presc_rst <= reset_presc;
	
	presc_in_buf : BUFG
               port map
                (O   => presc_in,
                 I   => presc_in_unbuffered);
	
	presc_inst : entity work.prescaler
		port map(clk_input  => presc_in,
			     clk_output => presc_out,
			     reset      => presc_rst,
			     presc      => presc_val);
	
	
	
	------------- BUFG -----------------
	--clock_out <= presc_out;
	
	clkout1_buf : BUFG
           port map
            (O   => clock_out,
             I   => presc_out);

end architecture RTL;
